[Font]
Font=
Name=Courier New
Size=9

[Assembler]
Assembler=
ForeGround=$00ff00
BackGround=$800000

[Comment]
Comment=
ForeGround=$c0c0c0
BackGround=$800000

[Directive]
Directive=
ForeGround=$ffffff
BackGround=$800000

[Identifier]
Identifier=
ForeGround=$00ffff
BackGround=$800000

[Invalid]
Invalid=
ForeGround=$ffffff
BackGround=$0000FF

[Key]
Key=
ForeGround=$ffffff
BackGround=$800000

[Number]
Number=
ForeGround=$00ffff
BackGround=$800000

[Space]
Space=
ForeGround=$800000
BackGround=$800000

[String]
String=
ForeGround=$00ffff
BackGround=$800000

[Symbol]
Symbol=
ForeGround=$ffffff
BackGround=$800000

[Editor]
Editor=
ForeGround=$80000005
BackGround=$800000
