[Font]
Name=Courier New
Size=9

[Assembler]
ForeGround=0
BackGround=$FFFFFF

[Comment]
ForeGround=0
BackGround=$FFFFFF

[Directive]
ForeGround=0
BackGround=$FFFFFF

[Identifier]
ForeGround=0
BackGround=$FFFFFF

[Invalid]
ForeGround=0
BackGround=$FFFFFF

[Key]
ForeGround=0
BackGround=$FFFFFF

[Number]
ForeGround=0
BackGround=$FFFFFF

[Space]
ForeGround=0
BackGround=$FFFFFF

[String]
ForeGround=0
BackGround=$FFFFFF

[Symbol]
ForeGround=0
BackGround=$FFFFFF

[Editor]
ForeGround=$000000
BackGround=$FFFFFF