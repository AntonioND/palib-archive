[Font]
Font=
Name=Courier New
Size=9

[Assembler]
Assembler=
ForeGround=$ff0000
BackGround=$ffff00

[Comment]
Comment=
ForeGround=$808080
BackGround=$ffff00

[Directive]
Directive=
ForeGround=$000000
BackGround=$ffff00

[Identifier]
Identifier=
ForeGround=$ff0000
BackGround=$ffff00

[Invalid]
Invalid=
ForeGround=$ffffff
BackGround=$0000FF

[Key]
Key=
ForeGround=$000000
BackGround=$ffff00

[Number]
Number=
ForeGround=$008080
BackGround=$ffff00

[Space]
Space=
ForeGround=$ffff00
BackGround=$ffff00

[String]
String=
ForeGround=$800080
BackGround=$ffff00

[Symbol]
Symbol=
ForeGround=$ff0000
BackGround=$ffff00

[Editor]
Editor=
ForeGround=$000000
BackGround=$ffff00
